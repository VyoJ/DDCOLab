module buffergate (y,a);  
input a;
output y;
assign y = a;
endmodule